------------------------------------------------------------------------------------------------------------
-- File name   : ucat_tb.vhd
--
-- Project     : EELE367 - Logic Design
--               uCat Final Project
--
-- Description : ModelSim test bench for ucat.vhd
--
-- Author(s)   : 	Matthew Handley
--
-- Note(s)     : 
--               
--
------------------------------------------------------------------------------------------------------------

entity ucat_tb is
end entity;

architecture ucat_tb_arch of ucat_tb is
  
  begin
    
    
    
end architecture;